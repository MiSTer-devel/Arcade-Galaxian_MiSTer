library ieee;
use ieee.std_logic_1164.all;

package sine_package is

	subtype table_value_type is integer range 0 to 16383;
	subtype table_index_type is std_logic_vector( 6 downto 0 );

	function get_table_value (table_index: table_index_type) return table_value_type;

end;

package body sine_package is

	function get_table_value (table_index: table_index_type) return table_value_type is
		variable table_value: table_value_type;
	begin
		case table_index is
			when "0000000" =>	table_value := 101;
			when "0000001" =>	table_value := 302;
			when "0000010" =>	table_value := 503;
			when "0000011" =>	table_value := 703;
			when "0000100" =>	table_value := 904;
			when "0000101" =>	table_value := 1105;
			when "0000110" =>	table_value := 1305;
			when "0000111" =>	table_value := 1506;
			when "0001000" =>	table_value := 1706;
			when "0001001" =>	table_value := 1906;
			when "0001010" =>	table_value := 2105;
			when "0001011" =>	table_value := 2304;
			when "0001100" =>	table_value := 2503;
			when "0001101" =>	table_value := 2702;
			when "0001110" =>	table_value := 2900;
			when "0001111" =>	table_value := 3098;
			when "0010000" =>	table_value := 3295;
			when "0010001" =>	table_value := 3491;
			when "0010010" =>	table_value := 3688;
			when "0010011" =>	table_value := 3883;
			when "0010100" =>	table_value := 4078;
			when "0010101" =>	table_value := 4273;
			when "0010110" =>	table_value := 4466;
			when "0010111" =>	table_value := 4659;
			when "0011000" =>	table_value := 4852;
			when "0011001" =>	table_value := 5044;
			when "0011010" =>	table_value := 5234;
			when "0011011" =>	table_value := 5425;
			when "0011100" =>	table_value := 5614;
			when "0011101" =>	table_value := 5802;
			when "0011110" =>	table_value := 5990;
			when "0011111" =>	table_value := 6177;
			when "0100000" =>	table_value := 6362;
			when "0100001" =>	table_value := 6547;
			when "0100010" =>	table_value := 6731;
			when "0100011" =>	table_value := 6914;
			when "0100100" =>	table_value := 7095;
			when "0100101" =>	table_value := 7276;
			when "0100110" =>	table_value := 7456;
			when "0100111" =>	table_value := 7634;
			when "0101000" =>	table_value := 7811;
			when "0101001" =>	table_value := 7988;
			when "0101010" =>	table_value := 8162;
			when "0101011" =>	table_value := 8336;
			when "0101100" =>	table_value := 8509;
			when "0101101" =>	table_value := 8680;
			when "0101110" =>	table_value := 8850;
			when "0101111" =>	table_value := 9018;
			when "0110000" =>	table_value := 9185;
			when "0110001" =>	table_value := 9351;
			when "0110010" =>	table_value := 9515;
			when "0110011" =>	table_value := 9678;
			when "0110100" =>	table_value := 9840;
			when "0110101" =>	table_value := 10000;
			when "0110110" =>	table_value := 10158;
			when "0110111" =>	table_value := 10315;
			when "0111000" =>	table_value := 10471;
			when "0111001" =>	table_value := 10625;
			when "0111010" =>	table_value := 10777;
			when "0111011" =>	table_value := 10927;
			when "0111100" =>	table_value := 11076;
			when "0111101" =>	table_value := 11224;
			when "0111110" =>	table_value := 11369;
			when "0111111" =>	table_value := 11513;
			when "1000000" =>	table_value := 11655;
			when "1000001" =>	table_value := 11796;
			when "1000010" =>	table_value := 11934;
			when "1000011" =>	table_value := 12071;
			when "1000100" =>	table_value := 12206;
			when "1000101" =>	table_value := 12339;
			when "1000110" =>	table_value := 12471;
			when "1000111" =>	table_value := 12600;
			when "1001000" =>	table_value := 12728;
			when "1001001" =>	table_value := 12853;
			when "1001010" =>	table_value := 12977;
			when "1001011" =>	table_value := 13099;
			when "1001100" =>	table_value := 13219;
			when "1001101" =>	table_value := 13336;
			when "1001110" =>	table_value := 13452;
			when "1001111" =>	table_value := 13566;
			when "1010000" =>	table_value := 13678;
			when "1010001" =>	table_value := 13787;
			when "1010010" =>	table_value := 13895;
			when "1010011" =>	table_value := 14000;
			when "1010100" =>	table_value := 14104;
			when "1010101" =>	table_value := 14205;
			when "1010110" =>	table_value := 14304;
			when "1010111" =>	table_value := 14401;
			when "1011000" =>	table_value := 14496;
			when "1011001" =>	table_value := 14588;
			when "1011010" =>	table_value := 14679;
			when "1011011" =>	table_value := 14767;
			when "1011100" =>	table_value := 14853;
			when "1011101" =>	table_value := 14936;
			when "1011110" =>	table_value := 15018;
			when "1011111" =>	table_value := 15097;
			when "1100000" =>	table_value := 15174;
			when "1100001" =>	table_value := 15249;
			when "1100010" =>	table_value := 15321;
			when "1100011" =>	table_value := 15391;
			when "1100100" =>	table_value := 15459;
			when "1100101" =>	table_value := 15524;
			when "1100110" =>	table_value := 15587;
			when "1100111" =>	table_value := 15648;
			when "1101000" =>	table_value := 15706;
			when "1101001" =>	table_value := 15762;
			when "1101010" =>	table_value := 15816;
			when "1101011" =>	table_value := 15867;
			when "1101100" =>	table_value := 15916;
			when "1101101" =>	table_value := 15963;
			when "1101110" =>	table_value := 16007;
			when "1101111" =>	table_value := 16048;
			when "1110000" =>	table_value := 16088;
			when "1110001" =>	table_value := 16124;
			when "1110010" =>	table_value := 16159;
			when "1110011" =>	table_value := 16191;
			when "1110100" =>	table_value := 16220;
			when "1110101" =>	table_value := 16247;
			when "1110110" =>	table_value := 16272;
			when "1110111" =>	table_value := 16294;
			when "1111000" =>	table_value := 16314;
			when "1111001" =>	table_value := 16331;
			when "1111010" =>	table_value := 16346;
			when "1111011" =>	table_value := 16358;
			when "1111100" =>	table_value := 16368;
			when "1111101" =>	table_value := 16375;
			when "1111110" =>	table_value := 16380;
			when "1111111" =>	table_value := 16383;
			when others => null;
		end case;
		return table_value;
	end;

end;
